library ieee;
use ieee.std_logic_1164.all;
entity store is
port (state: in std_logic_vector(2 downto 0);  --���뵱ǰ���״̬
	  s1,s2,s3,s4,s5,s6,s7,s8: out std_logic_vector(7 downto 0));  --���ҵ���Ӧ��ĸ�ĵ�����Ϣ�����
end store;

architecture behave of store is
begin

process(state)
begin
case state is
	when "001" =>   s1<="01000010";--������ʾH
					s2<="01000010";
					s3<="01000010";
					s4<="01000010";
					s5<="01111110";
					s6<="01000010";
					s7<="01000010";
					s8<="01000010";
	when "010" =>   s1<="00110000";--������ʾJ
					s2<="01001000";
					s3<="00001000";
					s4<="00001000";
					s5<="00001000";
					s6<="00001000";
					s7<="00001000";
					s8<="01111111";
	when "011" =>   s1<="01111100";--������ʾB
					s2<="01000010";
					s3<="01000010";
					s4<="01000100";
					s5<="01111000";
					s6<="01000100";
					s7<="01000100";
					s8<="01111000";
	when "100" =>   s1<="00001000";--������ʾT
					s2<="00001000";
					s3<="00001000";
					s4<="00001000";
					s5<="00001000";
					s6<="00001000";
					s7<="00001000";
					s8<="01111111";
	when "101" =>   s1<="11111111";--������ʾZ
					s2<="01000000";
					s3<="00100000";
					s4<="00010000";
					s5<="00001000";
					s6<="00000100";
					s7<="00000010";
					s8<="11111111";
	when others=>   s1<="00000000";--������ʾ
					s2<="00000000";
					s3<="00000000";
					s4<="00000000";
					s5<="00000000";
					s6<="00000000";
					s7<="00000000";
					s8<="00000000";
end case;
end process;

end behave;